`timescale 1ns / 1ns

module test(input logic a, b, output logic o);
    assign o = a ^ b;
endmodule